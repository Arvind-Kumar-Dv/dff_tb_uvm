typedef uvm_sequencer#(dff_tb_tx) dff_tb_sqr;
